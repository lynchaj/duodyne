-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

library ieee;
use ieee.std_logic_1164.all;
library altera;
use altera.altera_syn_attributes.all;

entity First is
	port
	(
-- {ALTERA_IO_BEGIN} DO NOT REMOVE THIS LINE!

		CK : out std_logic;
		CKDiv2 : out std_logic;
		CKDiv4 : out std_logic;
		CKDiv8 : out std_logic;
		CKDiv16 : out std_logic;
		Clock : in std_logic;
		Output_0 : out std_logic;
		Output_1 : out std_logic;
		Output_2 : out std_logic;
		Output_3 : out std_logic;
		Output_4 : out std_logic;
		Output_5 : out std_logic;
		Output_6 : out std_logic;
		Output_7 : out std_logic;
		Output_8 : out std_logic;
		Output_9 : out std_logic;
		Output_10 : out std_logic;
		Output_11 : out std_logic;
		Output_12 : out std_logic;
		Output_13 : out std_logic;
		Output_14 : out std_logic;
		Output_15 : out std_logic;
		Output_16 : out std_logic;
		Output_17 : out std_logic;
		Output_18 : out std_logic;
		Output_19 : out std_logic;
		Output_20 : out std_logic;
		Output_21 : out std_logic;
		Output_22 : out std_logic;
		Output_23 : out std_logic;
		Output_24 : out std_logic;
		Output_25 : out std_logic;
		Output_26 : out std_logic;
		Output_27 : out std_logic;
		Output_28 : out std_logic;
		Output_29 : out std_logic;
		Output_30 : out std_logic;
		Output_31 : out std_logic;
		Output_32 : out std_logic;
		Output_33 : out std_logic;
		Output_34 : out std_logic;
		Output_35 : out std_logic;
		Output_36 : out std_logic;
		Output_37 : out std_logic;
		Switch_1_0 : in std_logic;
		Switch_1_1 : in std_logic;
		Switch_1_2 : in std_logic;
		Switch_1_3 : in std_logic;
		Switch_1_4 : in std_logic;
		Switch_1_5 : in std_logic;
		Switch_1_6 : in std_logic;
		Switch_1_7 : in std_logic;
		Switch_2_0 : in std_logic;
		Switch_2_1 : in std_logic;
		Switch_2_2 : in std_logic;
		Switch_2_3 : in std_logic;
		Switch_2_4 : in std_logic;
		Switch_2_5 : in std_logic;
		Switch_2_6 : in std_logic;
		Switch_2_7 : in std_logic;
		TCK : in std_logic;
		TDI : in std_logic;
		TDO : out std_logic;
		TMS : in std_logic
-- {ALTERA_IO_END} DO NOT REMOVE THIS LINE!

	);

-- {ALTERA_ATTRIBUTE_BEGIN} DO NOT REMOVE THIS LINE!
-- {ALTERA_ATTRIBUTE_END} DO NOT REMOVE THIS LINE!
end First;

architecture ppl_type of First is

-- {ALTERA_COMPONENTS_BEGIN} DO NOT REMOVE THIS LINE!
-- {ALTERA_COMPONENTS_END} DO NOT REMOVE THIS LINE!
begin
-- {ALTERA_INSTANTIATION_BEGIN} DO NOT REMOVE THIS LINE!
-- {ALTERA_INSTANTIATION_END} DO NOT REMOVE THIS LINE!

end;
