library verilog;
use verilog.vl_types.all;
entity First_vlg_vec_tst is
end First_vlg_vec_tst;
